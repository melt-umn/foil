grammar edu:umn:cs:melt:foil:host:silverconstruction;

imports silver:langutil;
imports silver:langutil:pp;
imports silver:reflect;

imports silver:compiler:metatranslation;

imports silver:compiler:definition:core as silver;
imports silver:compiler:extension:patternmatching as silver;
imports edu:umn:cs:melt:foil:host:concretesyntax as foil;
imports edu:umn:cs:melt:foil:host:common as com;
imports edu:umn:cs:melt:foil:host:langs:ext as ext;
imports edu:umn:cs:melt:foil:host:langs:core as core;
