grammar edu:umn:cs:melt:foil:host:passes:ctrans;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:foil:host:common;
imports edu:umn:cs:melt:foil:host:langs:l1 as l1;
imports edu:umn:cs:melt:foil:host:langs:l2;
imports edu:umn:cs:melt:foil:host:passes:toL2;

synthesized attribute translation::Document;
synthesized attribute translations::[Document];
