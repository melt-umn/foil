grammar edu:umn:cs:melt:foil:host;

imports edu:umn:cs:melt:foil:host:langs:core;
imports edu:umn:cs:melt:foil:host:langs:ext;
imports edu:umn:cs:melt:foil:host:driver;

-- Export so that we can directly include this grammar in a parser
exports edu:umn:cs:melt:foil:host:concretesyntax;
