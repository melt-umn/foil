grammar edu:umn:cs:melt:foil:host:common;

imports silver:util:treemap as tm;
imports silver:langutil;
imports silver:langutil:pp;

-- This grammar contains common utilities that are shared across languages.
