grammar edu:umn:cs:melt:foil:extensions:records;
