grammar edu:umn:cs:melt:foil:host:concretesyntax;

imports edu:umn:cs:melt:foil:host:common as com;
imports edu:umn:cs:melt:foil:host:langs:ext as ext;

imports silver:langutil;
imports silver:langutil:lsp as lsp;
