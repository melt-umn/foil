grammar edu:umn:cs:melt:foil:host:concretesyntax;

