grammar edu:umn:cs:melt:foil:host:abstractsyntax:core;

tracked nonterminal Expr with pp, env, type, errors;
propagate errors on Expr;
