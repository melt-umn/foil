grammar edu:umn:cs:melt:foil:host:driver;

