grammar edu:umn:cs:melt:foil:host:langs:core;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:foil:host:common;
