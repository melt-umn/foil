grammar edu:umn:cs:melt:foil:host:abstractsyntax:core;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:foil:host:env;

