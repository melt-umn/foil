grammar edu:umn:cs:melt:foil:host:abstractsyntax:core;

tracked nonterminal Expr with pp, env, type, errors;
propagate env on Expr excluding let_;
propagate errors on Expr;

production var
top::Expr ::= n::Name
{
  top.pp = n.pp;
  top.type = n.lookupValue.type;
  top.errors <- n.lookupValue.lookupErrors;
}
production let_
top::Expr ::= d::VarDecl b::Expr
{
  top.pp = pp"let${groupnestlines(2, d.pp)}in${groupnestlines(2, b.pp)}end";
  top.type = b.type;
  d.env = top.env;
  b.env = addEnv(d.defs, top.env);
}

-- Literals
production intLit
top::Expr ::= i::Integer
{
  top.pp = pp"${i}";
  top.type = intType();
}
production floatLit
top::Expr ::= f::Float
{
  top.pp = pp"${f}";
  top.type = floatType();
}
production trueLit
top::Expr ::=
{
  top.pp = pp"true";
  top.type = boolType();
}
production falseLit
top::Expr ::=
{
  top.pp = pp"false";
  top.type = boolType();
}
production stringLit
top::Expr ::= s::String
{
  top.pp = pp"${s}";
  top.type = stringType();
}

-- Operators
production intAddOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) + (${e2})";
  top.type = intType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"+ expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"+ expected an int operand, but got ${show(80, e2.type)}")];
}
production intSubOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) - (${e2})";
  top.type = intType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"- expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"- expected an int operand, but got ${show(80, e2.type)}")];
}
production intMulOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) * (${e2})";
  top.type = intType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"* expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"* expected an int operand, but got ${show(80, e2.type)}")];
}
production intDivOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) / (${e2})";
  top.type = intType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"/ expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"/ expected an int operand, but got ${show(80, e2.type)}")];
}
production intEqOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) == (${e2})";
  top.type = boolType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"== expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"== expected an int operand, but got ${show(80, e2.type)}")];
}
production intNeqOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) != (${e2})";
  top.type = boolType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"!= expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"!= expected an int operand, but got ${show(80, e2.type)}")];
}
production intGtOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) > (${e2})";
  top.type = boolType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"> expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"> expected an int operand, but got ${show(80, e2.type)}")];
}
production intLtOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) < (${e2})";
  top.type = boolType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"< expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"< expected an int operand, but got ${show(80, e2.type)}")];
}
production intGteOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) >= (${e2})";
  top.type = boolType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s">= expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s">= expected an int operand, but got ${show(80, e2.type)}")];
}
production intLteOp
top::Expr ::= e1::Expr e2::Expr
{
  top.pp = pp"(${e1}) <= (${e2})";
  top.type = boolType();
  top.errors <-
    if e1.type == intType() then []
    else [errFromOrigin(e1, s"<= expected an int operand, but got ${show(80, e1.type)}")];
  top.errors <-
    if e2.type == intType() then []
    else [errFromOrigin(e2, s"<= expected an int operand, but got ${show(80, e2.type)}")];
}
