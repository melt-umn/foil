grammar edu:umn:cs:melt:foil:extensions:records;

imports edu:umn:cs:melt:foil:host:concretesyntax as cnc;
imports edu:umn:cs:melt:foil:host:langs:ext;
imports edu:umn:cs:melt:foil:host:langs:core as core;

imports silver:langutil;
imports silver:langutil:pp;
